`define EXP_OVERFLOW    1
`define EXP_DIVZERO     2 
`define EXP_BREAK       3
`define EXP_SYSCALL     4
`define EXP_ADDRERR     5
`define EXP_ERET        6
`define EXP_NOP         7
`define EXP_RESERVED    8

`define ALU_NOP         0
`define ALU_ADD         1
`define ALU_ADDI        2
`define ALU_ADDU        3
`define ALU_ADDIU       4
`define ALU_SUB         5
`define ALU_SUBU        6
`define ALU_SLT         7
`define ALU_SLTI        8
`define ALU_SLTU        9
`define ALU_SLTIU       10
`define ALU_DIV         11
`define ALU_DIVU        12
`define ALU_MULT        13
`define ALU_MULTU       14
`define ALU_AND         15
`define ALU_ANDI        16
`define ALU_LUI         17
`define ALU_NOR         18
`define ALU_OR          19
`define ALU_ORI         20
`define ALU_XOR         21
`define ALU_XORI        22
`define ALU_SLL         23
`define ALU_SLLV        24
`define ALU_SRA         25
`define ALU_SRAV        26
`define ALU_SRL         27
`define ALU_SRLV        28
`define ALU_BEQ         29
`define ALU_BNE         30
`define ALU_BGEZ        31
`define ALU_BGTZ        32
`define ALU_BLEZ        33
`define ALU_BLTZ        34
`define ALU_BLTZAL      35
`define ALU_BGEZAL      36
`define ALU_J           37
`define ALU_JAL         38
`define ALU_JR          39
`define ALU_JALR        40 
`define ALU_MFHI        41
`define ALU_MFLO        42
`define ALU_MTHI        43
`define ALU_MTLO        44
`define ALU_BREAK       45
`define ALU_SYSCALL     46
`define ALU_LB          47
`define ALU_LBU         48
`define ALU_LH          49
`define ALU_LHU         50
`define ALU_LW          51
`define ALU_SB          52
`define ALU_SH          53
`define ALU_SW          54
`define ALU_ERET        55
`define ALU_MFC0        56
`define ALU_MTC0        57
`define ALU_MUL         58

