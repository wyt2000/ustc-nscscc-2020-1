`define CLEAN_ALL_1 7
`define CLEAN_ALL_2 6
`define STALL_ALL   5
`define STALL_MEM   4
`define STALL_EX    3
`define STALL_ID    2
`define STALL_IF    1
`define STALL_IDLE  0

